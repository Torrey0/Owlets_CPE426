//Nothing to sim yet
